library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity op_block is
port (
	clock : in STD_LOGIC
	
	);
end op_block;

architecture Behavioral of op_block is

	

begin

	
	
end Behavioral;

